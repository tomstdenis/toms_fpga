//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 Education
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Sat Feb 14 11:31:51 2026

module Gowin_DPB (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [7:0] douta;
output [7:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [11:0] ada;
input [7:0] dina;
input [11:0] adb;
input [7:0] dinb;

wire [11:0] dpb_inst_0_douta_w;
wire [11:0] dpb_inst_0_doutb_w;
wire [11:0] dpb_inst_1_douta_w;
wire [11:0] dpb_inst_1_doutb_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[11:0],douta[3:0]}),
    .DOB({dpb_inst_0_doutb_w[11:0],doutb[3:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3:0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b0;
defparam dpb_inst_0.READ_MODE1 = 1'b0;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 4;
defparam dpb_inst_0.BIT_WIDTH_1 = 4;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h01110212FA01311F201B28050C0111E01FF0F720F10BAAE0998131D0B9A11006;
defparam dpb_inst_0.INIT_RAM_01 = 256'h6666666666666666666666660ADE5DF3C570AD14C2F70FCC580D0E1A90180DF2;
defparam dpb_inst_0.INIT_RAM_02 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_03 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_04 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_05 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_06 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_07 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_08 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_09 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_0A = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_0B = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_0C = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_0D = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_0E = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_0F = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_10 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_11 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_12 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_13 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_14 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_15 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_16 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_17 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_18 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_19 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_1A = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_1B = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_1C = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_1D = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_1E = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_1F = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_20 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_21 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_22 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_23 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_24 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_25 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_26 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_27 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_28 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_29 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_2A = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_2B = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_2C = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_2D = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_2E = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_2F = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_30 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_31 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_32 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_33 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_34 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_35 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_36 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_37 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_38 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_39 = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_3A = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_3B = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_3C = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_3D = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_3E = 256'h6666666666666666666666666666666666666666666666666666666666666666;
defparam dpb_inst_0.INIT_RAM_3F = 256'h6666666666666666666666666666666666666666666666666666666666666666;

DPB dpb_inst_1 (
    .DOA({dpb_inst_1_douta_w[11:0],douta[7:4]}),
    .DOB({dpb_inst_1_doutb_w[11:0],doutb[7:4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:4]})
);

defparam dpb_inst_1.READ_MODE0 = 1'b0;
defparam dpb_inst_1.READ_MODE1 = 1'b0;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 4;
defparam dpb_inst_1.BIT_WIDTH_1 = 4;
defparam dpb_inst_1.BLK_SEL_0 = 3'b000;
defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'h8E23D190EC819E0EE8E91080A1D1901D9EF8F84B8008488084808180848E0808;
defparam dpb_inst_1.INIT_RAM_01 = 256'hEEEEEEEEEEEEEEEEEEEEEEEE0002666666500024454524444405040E2A14C8EE;
defparam dpb_inst_1.INIT_RAM_02 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_03 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_04 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_05 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_06 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_07 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_08 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_09 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_0A = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_0B = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_0C = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_0D = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_0E = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_0F = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_10 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_11 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_12 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_13 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_14 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_15 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_16 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_17 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_18 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_19 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_1A = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_1B = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_1C = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_1D = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_1E = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_1F = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_20 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_21 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_22 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_23 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_24 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_25 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_26 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_27 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_28 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_29 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_2A = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_2B = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_2C = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_2D = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_2E = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_2F = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_30 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_31 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_32 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_33 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_34 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_35 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_36 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_37 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_38 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_39 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_3A = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_3B = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_3C = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_3D = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_3E = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam dpb_inst_1.INIT_RAM_3F = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;

endmodule //Gowin_DPB
