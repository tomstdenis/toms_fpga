module top(
    input clk,
    input rx_pin,
    output tx_pin,
    output led
);


endmodule