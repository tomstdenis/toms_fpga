`timescale 1ns/1ps

module useq_tb();


// Memory storage
    reg [7:0] mem [0:4095];
    
    // Latched data registers to simulate the 1-cycle BRAM latency
    reg [7:0] douta_reg;
    reg [7:0] doutb_reg;

    // The CPU sees the latched data
    wire [15:0] mem_data = {doutb_reg, douta_reg};
	wire wren;
	wire [7:0]  mem_out;
	wire [11:0] mem_addr;
	wire [11:0] mem_addr_next;
	
	reg clk;
	reg rst_n;
	reg [7:0] i_port;
	wire [7:0] o_port;
	reg read_fifo;
	reg write_fifo;
	wire fifo_empty;
	wire fifo_full;
	wire [7:0] fifo_out;
	reg [7:0] fifo_in;
	wire o_port_pulse;

    // Synchronous memory read: mimics Gowin DPB in Normal/Bypass mode
    always @(posedge clk) begin
        if (!rst_n) begin
            douta_reg <= 8'h00;
            doutb_reg <= 8'h00;
        end else begin
			// The memory array is sampled on the posedge
			if (wren) begin
				mem[mem_addr] <= mem_out;
			end else begin
				// Data becomes available for the CPU at the NEXT posedge
				douta_reg <= mem[mem_addr];
				doutb_reg <= mem[mem_addr_next]; // portB only reads if !wren to avoid SRAM address conflicts (can't read from address you're writing to)
			end
        end
    end

	useq #(.FIFO_DEPTH(16), .STACK_DEPTH(16), .ISR_VECT(12'hFE0), .ENABLE_IRQ(1), .ENABLE_HOST_FIFO_CTRL(1)) useq_dut(
		.clk(clk), .rst_n(rst_n), 
		.mem_data(mem_data), .i_port(i_port), 
		.mem_addr(mem_addr), .wren(wren), .mem_out(mem_out), .mem_addr_next(mem_addr_next), .o_port(o_port), .o_port_pulse(o_port_pulse),
		.read_fifo(read_fifo), .write_fifo(write_fifo), .fifo_empty(fifo_empty), .fifo_full(fifo_full),
		.fifo_out(fifo_out), .fifo_in(fifo_in));

    // Parameters for the simulation
    localparam CLK_PERIOD = 20; // 50MHz Clock
    // Clock Generation
    always #(CLK_PERIOD/2) clk = ~clk;

    // --- Verification Logic ---
    reg [9:0] T_PC;
    reg [7:0] T_A;
    reg [7:0] T_LR;
    reg [7:0] T_ILR;
    reg [7:0] T_R [15:0];
    
	integer i;
	integer j;
    initial begin
        // Setup for OSS CAD (GTKWave)
        $dumpfile("useq.vcd");
        $dumpvars(0, useq_tb);
		i_port = 0;
/*
		$readmemh("test1_clean.hex", mem);
		i_port = 8'hAB;
		reset_cpu();
		repeat(48) step_cpu();
		
		$display("Trying out interrupts...");
		$readmemh("test2_clean.hex", mem);
		i_port = 8'h00;
		reset_cpu();
		repeat(10) step_cpu();
		$display("Should be triggering an IRQ now...\n");
		i_port = 8'h01;
		repeat(20) step_cpu(); // ensure IRQ doesn't trip again
		$display("Should be triggering another IRQ now...\n");
		i_port = 8'h02;
		repeat(20) step_cpu(); // ensure IRQ doesn't trip again
		$display("Should be triggering last IRQ now (back on pin 0)...\n");
		i_port = 8'h01;
		repeat(20) step_cpu(); // ensure IRQ doesn't trip again
		$display("Should NOT be triggering last IRQ now (on pin 7)...\n");
		i_port = 8'h80;
		repeat(20) step_cpu(); // ensure IRQ doesn't trip again
        
		$display("Trying out FIFOS...");
		$readmemh("test3_clean.hex", mem);
		reset_cpu();
		step_cpu();
		write_fifo = 1;
		fifo_in = 8'hCC;
		step_cpu();
		write_fifo = 0;
		step_cpu();
		write_fifo = 1;
		fifo_in = 8'hDD;
		step_cpu();
		write_fifo = 0;
		repeat(16) step_cpu();
		read_fifo = 1;
		repeat(10) begin
			step_cpu();
			if (fifo_empty) read_fifo = 0;
		end
*/
		$display("Trying out uart demo...");
//		$readmemh("simple_clean.hex", mem);
		$readmemh("uart_clean.hex", mem);
		reset_cpu();
		repeat(131072) step_cpu();
		$finish;
	end

    task step_cpu();
		integer x;reg [11:0] ttpc;
		begin
			ttpc = useq_dut.PC;
			@(posedge clk);
			if (useq_dut.state == 2) begin
				$write("CPU: S=%d inst=%2h PC=%2h, A=%2h SP=%2d ILR=%2h IM=%2h IP=%2h OP=%2h FO=%2h FE=%d FF=%d R=[", useq_dut.state, useq_dut.instruct, useq_dut.PC, useq_dut.A, useq_dut.SP, useq_dut.ILR, useq_dut.int_mask, i_port, o_port, fifo_out, fifo_empty, fifo_full);
				for (x = 0; x < 16; x++) begin
					$write("%2h", useq_dut.R[x]);
					if (x < 15) begin
						$write(" ");
					end
				end
				$write("]\n");
			end
		end
	endtask

	task reset_cpu();
		integer x;
		begin
			// Initialize signals
			clk = 0;
			rst_n = 0;
			read_fifo = 0;
			write_fifo = 0;
			fifo_in = 0;
			T_PC = 0;
			T_A = 0;
			T_LR = 0;
			T_ILR = 0;
			for (x = 0; x < 16; x++) begin
				T_R[x] = 0;
			end
		
			// Reset
			repeat(5) @(posedge clk);
			rst_n = 1;
		end
	endtask
endmodule

