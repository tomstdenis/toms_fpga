//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 Education
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Mon Feb  9 23:42:30 2026

module Gowin_ROM16 (dout, ad);

output [7:0] dout;
input [7:0] ad;

wire [0:0] rom16_inst_0_dout;
wire [1:1] rom16_inst_1_dout;
wire [2:2] rom16_inst_2_dout;
wire [3:3] rom16_inst_3_dout;
wire [4:4] rom16_inst_4_dout;
wire [5:5] rom16_inst_5_dout;
wire [6:6] rom16_inst_6_dout;
wire [7:7] rom16_inst_7_dout;
wire [0:0] rom16_inst_8_dout;
wire [1:1] rom16_inst_9_dout;
wire [2:2] rom16_inst_10_dout;
wire [3:3] rom16_inst_11_dout;
wire [4:4] rom16_inst_12_dout;
wire [5:5] rom16_inst_13_dout;
wire [6:6] rom16_inst_14_dout;
wire [7:7] rom16_inst_15_dout;
wire [0:0] rom16_inst_16_dout;
wire [1:1] rom16_inst_17_dout;
wire [2:2] rom16_inst_18_dout;
wire [3:3] rom16_inst_19_dout;
wire [4:4] rom16_inst_20_dout;
wire [5:5] rom16_inst_21_dout;
wire [6:6] rom16_inst_22_dout;
wire [7:7] rom16_inst_23_dout;
wire [0:0] rom16_inst_24_dout;
wire [1:1] rom16_inst_25_dout;
wire [2:2] rom16_inst_26_dout;
wire [3:3] rom16_inst_27_dout;
wire [4:4] rom16_inst_28_dout;
wire [5:5] rom16_inst_29_dout;
wire [6:6] rom16_inst_30_dout;
wire [7:7] rom16_inst_31_dout;
wire [0:0] rom16_inst_32_dout;
wire [1:1] rom16_inst_33_dout;
wire [2:2] rom16_inst_34_dout;
wire [3:3] rom16_inst_35_dout;
wire [4:4] rom16_inst_36_dout;
wire [5:5] rom16_inst_37_dout;
wire [6:6] rom16_inst_38_dout;
wire [7:7] rom16_inst_39_dout;
wire [0:0] rom16_inst_40_dout;
wire [1:1] rom16_inst_41_dout;
wire [2:2] rom16_inst_42_dout;
wire [3:3] rom16_inst_43_dout;
wire [4:4] rom16_inst_44_dout;
wire [5:5] rom16_inst_45_dout;
wire [6:6] rom16_inst_46_dout;
wire [7:7] rom16_inst_47_dout;
wire [0:0] rom16_inst_48_dout;
wire [1:1] rom16_inst_49_dout;
wire [2:2] rom16_inst_50_dout;
wire [3:3] rom16_inst_51_dout;
wire [4:4] rom16_inst_52_dout;
wire [5:5] rom16_inst_53_dout;
wire [6:6] rom16_inst_54_dout;
wire [7:7] rom16_inst_55_dout;
wire [0:0] rom16_inst_56_dout;
wire [1:1] rom16_inst_57_dout;
wire [2:2] rom16_inst_58_dout;
wire [3:3] rom16_inst_59_dout;
wire [4:4] rom16_inst_60_dout;
wire [5:5] rom16_inst_61_dout;
wire [6:6] rom16_inst_62_dout;
wire [7:7] rom16_inst_63_dout;
wire [0:0] rom16_inst_64_dout;
wire [1:1] rom16_inst_65_dout;
wire [2:2] rom16_inst_66_dout;
wire [3:3] rom16_inst_67_dout;
wire [4:4] rom16_inst_68_dout;
wire [5:5] rom16_inst_69_dout;
wire [6:6] rom16_inst_70_dout;
wire [7:7] rom16_inst_71_dout;
wire [0:0] rom16_inst_72_dout;
wire [1:1] rom16_inst_73_dout;
wire [2:2] rom16_inst_74_dout;
wire [3:3] rom16_inst_75_dout;
wire [4:4] rom16_inst_76_dout;
wire [5:5] rom16_inst_77_dout;
wire [6:6] rom16_inst_78_dout;
wire [7:7] rom16_inst_79_dout;
wire [0:0] rom16_inst_80_dout;
wire [1:1] rom16_inst_81_dout;
wire [2:2] rom16_inst_82_dout;
wire [3:3] rom16_inst_83_dout;
wire [4:4] rom16_inst_84_dout;
wire [5:5] rom16_inst_85_dout;
wire [6:6] rom16_inst_86_dout;
wire [7:7] rom16_inst_87_dout;
wire [0:0] rom16_inst_88_dout;
wire [1:1] rom16_inst_89_dout;
wire [2:2] rom16_inst_90_dout;
wire [3:3] rom16_inst_91_dout;
wire [4:4] rom16_inst_92_dout;
wire [5:5] rom16_inst_93_dout;
wire [6:6] rom16_inst_94_dout;
wire [7:7] rom16_inst_95_dout;
wire [0:0] rom16_inst_96_dout;
wire [1:1] rom16_inst_97_dout;
wire [2:2] rom16_inst_98_dout;
wire [3:3] rom16_inst_99_dout;
wire [4:4] rom16_inst_100_dout;
wire [5:5] rom16_inst_101_dout;
wire [6:6] rom16_inst_102_dout;
wire [7:7] rom16_inst_103_dout;
wire [0:0] rom16_inst_104_dout;
wire [1:1] rom16_inst_105_dout;
wire [2:2] rom16_inst_106_dout;
wire [3:3] rom16_inst_107_dout;
wire [4:4] rom16_inst_108_dout;
wire [5:5] rom16_inst_109_dout;
wire [6:6] rom16_inst_110_dout;
wire [7:7] rom16_inst_111_dout;
wire [0:0] rom16_inst_112_dout;
wire [1:1] rom16_inst_113_dout;
wire [2:2] rom16_inst_114_dout;
wire [3:3] rom16_inst_115_dout;
wire [4:4] rom16_inst_116_dout;
wire [5:5] rom16_inst_117_dout;
wire [6:6] rom16_inst_118_dout;
wire [7:7] rom16_inst_119_dout;
wire [0:0] rom16_inst_120_dout;
wire [1:1] rom16_inst_121_dout;
wire [2:2] rom16_inst_122_dout;
wire [3:3] rom16_inst_123_dout;
wire [4:4] rom16_inst_124_dout;
wire [5:5] rom16_inst_125_dout;
wire [6:6] rom16_inst_126_dout;
wire [7:7] rom16_inst_127_dout;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;

ROM16 rom16_inst_0 (
    .DO(rom16_inst_0_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_0.INIT_0 = 16'hFFF3;

ROM16 rom16_inst_1 (
    .DO(rom16_inst_1_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_1.INIT_0 = 16'hFFEF;

ROM16 rom16_inst_2 (
    .DO(rom16_inst_2_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_2.INIT_0 = 16'hFFEB;

ROM16 rom16_inst_3 (
    .DO(rom16_inst_3_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_3.INIT_0 = 16'hFFEB;

ROM16 rom16_inst_4 (
    .DO(rom16_inst_4_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_4.INIT_0 = 16'h001D;

ROM16 rom16_inst_5 (
    .DO(rom16_inst_5_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_5.INIT_0 = 16'hFFE1;

ROM16 rom16_inst_6 (
    .DO(rom16_inst_6_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_6.INIT_0 = 16'h000E;

ROM16 rom16_inst_7 (
    .DO(rom16_inst_7_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_7.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_8 (
    .DO(rom16_inst_8_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_8.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_9 (
    .DO(rom16_inst_9_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_9.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_10 (
    .DO(rom16_inst_10_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_10.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_11 (
    .DO(rom16_inst_11_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_11.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_12 (
    .DO(rom16_inst_12_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_12.INIT_0 = 16'h0000;

ROM16 rom16_inst_13 (
    .DO(rom16_inst_13_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_13.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_14 (
    .DO(rom16_inst_14_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_14.INIT_0 = 16'h0000;

ROM16 rom16_inst_15 (
    .DO(rom16_inst_15_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_15.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_16 (
    .DO(rom16_inst_16_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_16.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_17 (
    .DO(rom16_inst_17_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_17.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_18 (
    .DO(rom16_inst_18_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_18.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_19 (
    .DO(rom16_inst_19_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_19.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_20 (
    .DO(rom16_inst_20_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_20.INIT_0 = 16'h0000;

ROM16 rom16_inst_21 (
    .DO(rom16_inst_21_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_21.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_22 (
    .DO(rom16_inst_22_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_22.INIT_0 = 16'h0000;

ROM16 rom16_inst_23 (
    .DO(rom16_inst_23_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_23.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_24 (
    .DO(rom16_inst_24_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_24.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_25 (
    .DO(rom16_inst_25_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_25.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_26 (
    .DO(rom16_inst_26_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_26.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_27 (
    .DO(rom16_inst_27_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_27.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_28 (
    .DO(rom16_inst_28_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_28.INIT_0 = 16'h0000;

ROM16 rom16_inst_29 (
    .DO(rom16_inst_29_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_29.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_30 (
    .DO(rom16_inst_30_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_30.INIT_0 = 16'h0000;

ROM16 rom16_inst_31 (
    .DO(rom16_inst_31_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_31.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_32 (
    .DO(rom16_inst_32_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_32.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_33 (
    .DO(rom16_inst_33_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_33.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_34 (
    .DO(rom16_inst_34_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_34.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_35 (
    .DO(rom16_inst_35_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_35.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_36 (
    .DO(rom16_inst_36_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_36.INIT_0 = 16'h0000;

ROM16 rom16_inst_37 (
    .DO(rom16_inst_37_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_37.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_38 (
    .DO(rom16_inst_38_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_38.INIT_0 = 16'h0000;

ROM16 rom16_inst_39 (
    .DO(rom16_inst_39_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_39.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_40 (
    .DO(rom16_inst_40_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_40.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_41 (
    .DO(rom16_inst_41_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_41.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_42 (
    .DO(rom16_inst_42_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_42.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_43 (
    .DO(rom16_inst_43_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_43.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_44 (
    .DO(rom16_inst_44_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_44.INIT_0 = 16'h0000;

ROM16 rom16_inst_45 (
    .DO(rom16_inst_45_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_45.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_46 (
    .DO(rom16_inst_46_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_46.INIT_0 = 16'h0000;

ROM16 rom16_inst_47 (
    .DO(rom16_inst_47_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_47.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_48 (
    .DO(rom16_inst_48_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_48.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_49 (
    .DO(rom16_inst_49_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_49.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_50 (
    .DO(rom16_inst_50_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_50.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_51 (
    .DO(rom16_inst_51_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_51.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_52 (
    .DO(rom16_inst_52_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_52.INIT_0 = 16'h0000;

ROM16 rom16_inst_53 (
    .DO(rom16_inst_53_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_53.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_54 (
    .DO(rom16_inst_54_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_54.INIT_0 = 16'h0000;

ROM16 rom16_inst_55 (
    .DO(rom16_inst_55_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_55.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_56 (
    .DO(rom16_inst_56_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_56.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_57 (
    .DO(rom16_inst_57_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_57.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_58 (
    .DO(rom16_inst_58_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_58.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_59 (
    .DO(rom16_inst_59_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_59.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_60 (
    .DO(rom16_inst_60_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_60.INIT_0 = 16'h0000;

ROM16 rom16_inst_61 (
    .DO(rom16_inst_61_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_61.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_62 (
    .DO(rom16_inst_62_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_62.INIT_0 = 16'h0000;

ROM16 rom16_inst_63 (
    .DO(rom16_inst_63_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_63.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_64 (
    .DO(rom16_inst_64_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_64.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_65 (
    .DO(rom16_inst_65_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_65.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_66 (
    .DO(rom16_inst_66_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_66.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_67 (
    .DO(rom16_inst_67_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_67.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_68 (
    .DO(rom16_inst_68_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_68.INIT_0 = 16'h0000;

ROM16 rom16_inst_69 (
    .DO(rom16_inst_69_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_69.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_70 (
    .DO(rom16_inst_70_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_70.INIT_0 = 16'h0000;

ROM16 rom16_inst_71 (
    .DO(rom16_inst_71_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_71.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_72 (
    .DO(rom16_inst_72_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_72.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_73 (
    .DO(rom16_inst_73_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_73.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_74 (
    .DO(rom16_inst_74_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_74.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_75 (
    .DO(rom16_inst_75_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_75.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_76 (
    .DO(rom16_inst_76_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_76.INIT_0 = 16'h0000;

ROM16 rom16_inst_77 (
    .DO(rom16_inst_77_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_77.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_78 (
    .DO(rom16_inst_78_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_78.INIT_0 = 16'h0000;

ROM16 rom16_inst_79 (
    .DO(rom16_inst_79_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_79.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_80 (
    .DO(rom16_inst_80_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_80.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_81 (
    .DO(rom16_inst_81_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_81.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_82 (
    .DO(rom16_inst_82_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_82.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_83 (
    .DO(rom16_inst_83_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_83.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_84 (
    .DO(rom16_inst_84_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_84.INIT_0 = 16'h0000;

ROM16 rom16_inst_85 (
    .DO(rom16_inst_85_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_85.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_86 (
    .DO(rom16_inst_86_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_86.INIT_0 = 16'h0000;

ROM16 rom16_inst_87 (
    .DO(rom16_inst_87_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_87.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_88 (
    .DO(rom16_inst_88_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_88.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_89 (
    .DO(rom16_inst_89_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_89.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_90 (
    .DO(rom16_inst_90_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_90.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_91 (
    .DO(rom16_inst_91_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_91.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_92 (
    .DO(rom16_inst_92_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_92.INIT_0 = 16'h0000;

ROM16 rom16_inst_93 (
    .DO(rom16_inst_93_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_93.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_94 (
    .DO(rom16_inst_94_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_94.INIT_0 = 16'h0000;

ROM16 rom16_inst_95 (
    .DO(rom16_inst_95_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_95.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_96 (
    .DO(rom16_inst_96_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_96.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_97 (
    .DO(rom16_inst_97_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_97.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_98 (
    .DO(rom16_inst_98_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_98.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_99 (
    .DO(rom16_inst_99_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_99.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_100 (
    .DO(rom16_inst_100_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_100.INIT_0 = 16'h0000;

ROM16 rom16_inst_101 (
    .DO(rom16_inst_101_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_101.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_102 (
    .DO(rom16_inst_102_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_102.INIT_0 = 16'h0000;

ROM16 rom16_inst_103 (
    .DO(rom16_inst_103_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_103.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_104 (
    .DO(rom16_inst_104_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_104.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_105 (
    .DO(rom16_inst_105_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_105.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_106 (
    .DO(rom16_inst_106_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_106.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_107 (
    .DO(rom16_inst_107_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_107.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_108 (
    .DO(rom16_inst_108_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_108.INIT_0 = 16'h0000;

ROM16 rom16_inst_109 (
    .DO(rom16_inst_109_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_109.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_110 (
    .DO(rom16_inst_110_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_110.INIT_0 = 16'h0000;

ROM16 rom16_inst_111 (
    .DO(rom16_inst_111_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_111.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_112 (
    .DO(rom16_inst_112_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_112.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_113 (
    .DO(rom16_inst_113_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_113.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_114 (
    .DO(rom16_inst_114_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_114.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_115 (
    .DO(rom16_inst_115_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_115.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_116 (
    .DO(rom16_inst_116_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_116.INIT_0 = 16'h0000;

ROM16 rom16_inst_117 (
    .DO(rom16_inst_117_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_117.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_118 (
    .DO(rom16_inst_118_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_118.INIT_0 = 16'h0000;

ROM16 rom16_inst_119 (
    .DO(rom16_inst_119_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_119.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_120 (
    .DO(rom16_inst_120_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_120.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_121 (
    .DO(rom16_inst_121_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_121.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_122 (
    .DO(rom16_inst_122_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_122.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_123 (
    .DO(rom16_inst_123_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_123.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_124 (
    .DO(rom16_inst_124_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_124.INIT_0 = 16'h0000;

ROM16 rom16_inst_125 (
    .DO(rom16_inst_125_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_125.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_126 (
    .DO(rom16_inst_126_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_126.INIT_0 = 16'h0000;

ROM16 rom16_inst_127 (
    .DO(rom16_inst_127_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_127.INIT_0 = 16'hFFFF;

MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(rom16_inst_0_dout[0]),
  .I1(rom16_inst_8_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(rom16_inst_16_dout[0]),
  .I1(rom16_inst_24_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(rom16_inst_32_dout[0]),
  .I1(rom16_inst_40_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(rom16_inst_48_dout[0]),
  .I1(rom16_inst_56_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(rom16_inst_64_dout[0]),
  .I1(rom16_inst_72_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(rom16_inst_80_dout[0]),
  .I1(rom16_inst_88_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(rom16_inst_96_dout[0]),
  .I1(rom16_inst_104_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(rom16_inst_112_dout[0]),
  .I1(rom16_inst_120_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(ad[5])
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(ad[5])
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(ad[5])
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(ad[5])
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(ad[6])
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(ad[6])
);
MUX2 mux_inst_14 (
  .O(dout[0]),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(ad[7])
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(rom16_inst_1_dout[1]),
  .I1(rom16_inst_9_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(rom16_inst_17_dout[1]),
  .I1(rom16_inst_25_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(rom16_inst_33_dout[1]),
  .I1(rom16_inst_41_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(rom16_inst_49_dout[1]),
  .I1(rom16_inst_57_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(rom16_inst_65_dout[1]),
  .I1(rom16_inst_73_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(rom16_inst_81_dout[1]),
  .I1(rom16_inst_89_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(rom16_inst_97_dout[1]),
  .I1(rom16_inst_105_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(rom16_inst_113_dout[1]),
  .I1(rom16_inst_121_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(mux_o_15),
  .I1(mux_o_16),
  .S0(ad[5])
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(mux_o_17),
  .I1(mux_o_18),
  .S0(ad[5])
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_19),
  .I1(mux_o_20),
  .S0(ad[5])
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_21),
  .I1(mux_o_22),
  .S0(ad[5])
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(mux_o_23),
  .I1(mux_o_24),
  .S0(ad[6])
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(mux_o_25),
  .I1(mux_o_26),
  .S0(ad[6])
);
MUX2 mux_inst_29 (
  .O(dout[1]),
  .I0(mux_o_27),
  .I1(mux_o_28),
  .S0(ad[7])
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(rom16_inst_2_dout[2]),
  .I1(rom16_inst_10_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(rom16_inst_18_dout[2]),
  .I1(rom16_inst_26_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(rom16_inst_34_dout[2]),
  .I1(rom16_inst_42_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(rom16_inst_50_dout[2]),
  .I1(rom16_inst_58_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(rom16_inst_66_dout[2]),
  .I1(rom16_inst_74_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(rom16_inst_82_dout[2]),
  .I1(rom16_inst_90_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(rom16_inst_98_dout[2]),
  .I1(rom16_inst_106_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(rom16_inst_114_dout[2]),
  .I1(rom16_inst_122_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(ad[5])
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(ad[5])
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_34),
  .I1(mux_o_35),
  .S0(ad[5])
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(mux_o_36),
  .I1(mux_o_37),
  .S0(ad[5])
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(ad[6])
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(ad[6])
);
MUX2 mux_inst_44 (
  .O(dout[2]),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(ad[7])
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(rom16_inst_3_dout[3]),
  .I1(rom16_inst_11_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(rom16_inst_19_dout[3]),
  .I1(rom16_inst_27_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(rom16_inst_35_dout[3]),
  .I1(rom16_inst_43_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(rom16_inst_51_dout[3]),
  .I1(rom16_inst_59_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(rom16_inst_67_dout[3]),
  .I1(rom16_inst_75_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(rom16_inst_83_dout[3]),
  .I1(rom16_inst_91_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(rom16_inst_99_dout[3]),
  .I1(rom16_inst_107_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(rom16_inst_115_dout[3]),
  .I1(rom16_inst_123_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(ad[5])
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_47),
  .I1(mux_o_48),
  .S0(ad[5])
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(ad[5])
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(ad[5])
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(mux_o_53),
  .I1(mux_o_54),
  .S0(ad[6])
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(mux_o_55),
  .I1(mux_o_56),
  .S0(ad[6])
);
MUX2 mux_inst_59 (
  .O(dout[3]),
  .I0(mux_o_57),
  .I1(mux_o_58),
  .S0(ad[7])
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(rom16_inst_4_dout[4]),
  .I1(rom16_inst_12_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(rom16_inst_20_dout[4]),
  .I1(rom16_inst_28_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(rom16_inst_36_dout[4]),
  .I1(rom16_inst_44_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(rom16_inst_52_dout[4]),
  .I1(rom16_inst_60_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(rom16_inst_68_dout[4]),
  .I1(rom16_inst_76_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(rom16_inst_84_dout[4]),
  .I1(rom16_inst_92_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(rom16_inst_100_dout[4]),
  .I1(rom16_inst_108_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(rom16_inst_116_dout[4]),
  .I1(rom16_inst_124_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(ad[5])
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(ad[5])
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(ad[5])
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(ad[5])
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(ad[6])
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(ad[6])
);
MUX2 mux_inst_74 (
  .O(dout[4]),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(ad[7])
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(rom16_inst_5_dout[5]),
  .I1(rom16_inst_13_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(rom16_inst_21_dout[5]),
  .I1(rom16_inst_29_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(rom16_inst_37_dout[5]),
  .I1(rom16_inst_45_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(rom16_inst_53_dout[5]),
  .I1(rom16_inst_61_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(rom16_inst_69_dout[5]),
  .I1(rom16_inst_77_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(rom16_inst_85_dout[5]),
  .I1(rom16_inst_93_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(rom16_inst_101_dout[5]),
  .I1(rom16_inst_109_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(rom16_inst_117_dout[5]),
  .I1(rom16_inst_125_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(mux_o_75),
  .I1(mux_o_76),
  .S0(ad[5])
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(ad[5])
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(ad[5])
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(ad[5])
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(ad[6])
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(ad[6])
);
MUX2 mux_inst_89 (
  .O(dout[5]),
  .I0(mux_o_87),
  .I1(mux_o_88),
  .S0(ad[7])
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(rom16_inst_6_dout[6]),
  .I1(rom16_inst_14_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(rom16_inst_22_dout[6]),
  .I1(rom16_inst_30_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(rom16_inst_38_dout[6]),
  .I1(rom16_inst_46_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(rom16_inst_54_dout[6]),
  .I1(rom16_inst_62_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(rom16_inst_70_dout[6]),
  .I1(rom16_inst_78_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(rom16_inst_86_dout[6]),
  .I1(rom16_inst_94_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(rom16_inst_102_dout[6]),
  .I1(rom16_inst_110_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(rom16_inst_118_dout[6]),
  .I1(rom16_inst_126_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(ad[5])
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(ad[5])
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(ad[5])
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_96),
  .I1(mux_o_97),
  .S0(ad[5])
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(ad[6])
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(ad[6])
);
MUX2 mux_inst_104 (
  .O(dout[6]),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(ad[7])
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(rom16_inst_7_dout[7]),
  .I1(rom16_inst_15_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(rom16_inst_23_dout[7]),
  .I1(rom16_inst_31_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(rom16_inst_39_dout[7]),
  .I1(rom16_inst_47_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(rom16_inst_55_dout[7]),
  .I1(rom16_inst_63_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(rom16_inst_71_dout[7]),
  .I1(rom16_inst_79_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(rom16_inst_87_dout[7]),
  .I1(rom16_inst_95_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(rom16_inst_103_dout[7]),
  .I1(rom16_inst_111_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(rom16_inst_119_dout[7]),
  .I1(rom16_inst_127_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(ad[5])
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(ad[5])
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(ad[5])
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_111),
  .I1(mux_o_112),
  .S0(ad[5])
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(ad[6])
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_115),
  .I1(mux_o_116),
  .S0(ad[6])
);
MUX2 mux_inst_119 (
  .O(dout[7]),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(ad[7])
);
endmodule //Gowin_ROM16
