module top(
    input clk,
    output pwm
);



endmodule