`timescale 1ns/1ps

module useq
#(parameter
	FIFO_DEPTH=16,
	ISR_VECT=12'hFE0,					// 32 bytes short of top of memory
	ENABLE_IRQ=1,
	ENABLE_HOST_FIFO_CTRL=1,
	STACK_DEPTH=16
)(
	input clk,
	input rst_n,
	
	input [15:0] mem_data,				// 16-bit input fed from {MEM[mem_addr_next}, MEM[mem_addr]}
	output reg wren,					// write enable on portA (uses mem_addr)
	output reg [7:0] mem_out,			// data to write to portA of memory
	input [7:0] i_port,					// input port you can connect other pins to feed data into the core

	input read_fifo,					// pulse this high to read a byte from the FIFO into fifo_out in the next clock cycle
	input write_fifo,					// pulse this high to write from fifo_in into the FIFO
	output fifo_empty,					// high when the FIFO is empty
	output fifo_full,					// high when the FIFO is full
	input [7:0] fifo_in,				// The FIFO input into the core when pulsing write_fifo 
	output reg [7:0] fifo_out,			// The fifo output from the core when pulsing read_fifo
	
	output reg [11:0] mem_addr,			// The address the core needs mem_data from in the next clock cycle
	output reg [11:0] mem_addr_next,
	output reg [7:0] o_port,			// output port you can connect other pins to feed data out of the core.
	output reg o_port_pulse				// This pin toggles when a write to o_port is done.
);

	reg [7:0] A;								// A accumulator
	reg [7:0] tA;								// temporaty A used for IRQ
	reg [7:0] tR[1:0];							// temporary R[0..1] used for IRQ
	reg [$clog2(STACK_DEPTH):0] SP;				// stack pointer
	reg [11:0] PC;								// PC program counter
	reg [8:0] T;								// T temporary register used for WAITA opcode
	reg [8:0] tT;								// copy of T for IRQ context switching
	reg [11:0] LR[STACK_DEPTH-1:0];				// LR link register
	reg [11:0] ILR;								// ILR IRQ link register
	reg [7:0] instruct;							// current opcode
	reg [7:0] instruct_imm;						// immediate for the instruction
	reg [7:0] R[15:0];							// R register file
	reg [7:0] l_i_port;							// latched copy of i_port
	reg [7:0] int_mask;							// The IRQ mask applied to i_port set by SEI opcode
	reg [11:0] isr_vect;						// Where to jump when an IRQ happens
	reg int_enable;								// Interrupt enable (set by SEI, disabled during IRQ)
	reg [7:0] FIFO[FIFO_DEPTH-1:0];				// Message passing FIFO
	reg [$clog2(FIFO_DEPTH)-1:0] fifo_rptr;		// FIFO read pointer
	reg [$clog2(FIFO_DEPTH)-1:0] fifo_wptr;		// FIFO write pointer
	reg [2:0] state;							// current FSM state

	localparam
		FETCH = 0,
		DECODE = 1,
		EXECUTE = 2,
		LOADA = 3,
		LOADA_REG = 4,
		STOREA = 5,
		LOADIND = 6,
		LOADIND_REG = 7;

	integer i;

	// exec1 wires
	wire [3:0] d_imm = instruct[3:0];
	wire [2:0] s_imm = instruct[3:1];
	wire       b_imm = instruct[0];

	wire		int_triggered = |((i_port & ~l_i_port) & int_mask) & int_enable & (ENABLE_IRQ ? 1'b1 : 1'b0);
	wire 		host_wants_fifo = read_fifo ^ write_fifo;
	assign		fifo_empty = (R[15] == 0) ? 1'b1 : 1'b0;
	assign		fifo_full = (R[15] == FIFO_DEPTH) ? 1'b1 : 1'b0;

	always @(posedge clk) begin
		if (!rst_n) begin
			if (ENABLE_IRQ == 1) begin
				tA <= 0;
				tR[0] <= 0;
				tR[1] <= 0;
				tT <= 0;
				ILR <= 0;
				int_mask <= 0;
				int_enable <= 0;
				isr_vect <= ISR_VECT;
			end
			A <= 0;
			PC <= 0;
			T <= 0;
			state <= FETCH;
			l_i_port <= 0;
			o_port <= 8'hff;
			instruct <= 8'hE6;
			instruct_imm <= 0;
			mem_addr <= 0;
			mem_addr_next <= 1;
			wren <= 0;
			o_port_pulse <= 0;
			for (i=0; i<16; i=i+1) begin
				R[i] <= 0;
			end
			for (i=0; i<FIFO_DEPTH; i=i+1) begin
				FIFO[i] <= 0;
			end
			SP <= 0;
			for (i=0; i<STACK_DEPTH; i=i+1) begin
				LR[i] <= 0;
			end
			fifo_rptr <= 0;
			fifo_wptr <= 0;
			fifo_out <= 0;
		end else begin
			if (ENABLE_HOST_FIFO_CTRL == 1 && host_wants_fifo) begin
				if (read_fifo) begin
					// read fifo to o_port
					if (R[15] != 0) begin
						fifo_out <= FIFO[fifo_rptr];
						fifo_rptr <= fifo_rptr + 1'b1;
						R[15] <= R[15] - 1'b1;
					end else begin
						// fifo empty so write 0 to the port
						o_port <= 8'd0;
					end
				end else begin
					if (R[15] != FIFO_DEPTH) begin
						FIFO[fifo_wptr] <= fifo_in;			// store fifo data
						fifo_wptr <= fifo_wptr + 1'b1;		// increment write pointer
						R[15] <= R[15] + 1'b1;				// increment fifo count
					end
				end
			end else begin
				l_i_port <= i_port;						// only latch port when we're running the CPU
				if (int_triggered) begin
					// we hit an interrupt, so disable further interrupts until an RTI
					int_enable <= 0;
					ILR <= PC;     			// save where we interrupted
					tA <= A;
					tR[0] <= R[0];
					tR[1] <= R[1];
					tT <= T;
					mem_addr <= isr_vect;	// jump to ISR vector
					mem_addr_next <= isr_vect + 12'd1;
					PC <= isr_vect;
					state <= FETCH;			// need another FETCH cycle
				end else begin
					case(state)
						FETCH:
							begin
								state <= DECODE;
							end							
						DECODE:
							begin
								instruct <= mem_data[7:0];
								instruct_imm <= mem_data[15:8];
								state <= EXECUTE;
							end
						EXECUTE:
							begin
								// no interrupt so jump here
								`include "exec1_top.v"
							end
						LOADA: // wait a cycle for the BRAM to respond
							begin
								state <= LOADA_REG;
							end
						LOADA_REG: // mem_addr was set to the address we want to load and store in A
							begin
								A <= mem_data[7:0];
								mem_addr <= PC;
								mem_addr_next <= PC + 12'd1;
								state <= FETCH;
							end
						STOREA: // Cycle after a store is initiated
							begin
								wren <= 0;
								mem_addr <= PC;
								mem_addr_next <= PC + 12'd1;
								state <= FETCH;
							end
						LOADIND:
							begin
								state <= LOADIND_REG;
							end
						LOADIND_REG: // load R14:R13 with memory and advance
							begin
								R[13] <= mem_data[7:0];
								R[14] <= mem_data[15:8];
								mem_addr <= PC;
								mem_addr_next <= PC + 12'd1;
								state <= FETCH;
							end
					endcase
				end
			end
		end
	end
endmodule

